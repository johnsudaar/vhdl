module hello_world ;

initial begin
  $display ( "Hello world by Johnsudaar" );
  #10 $finish;
end

endmodule
